magic
tech sky130B
magscale 1 2
timestamp 1697381458
<< obsli1 >>
rect 1104 2159 258888 137649
<< obsm1 >>
rect 934 1368 258888 137680
<< metal2 >>
rect 4434 139200 4490 140000
rect 8482 139200 8538 140000
rect 12530 139200 12586 140000
rect 16578 139200 16634 140000
rect 20626 139200 20682 140000
rect 24674 139200 24730 140000
rect 28722 139200 28778 140000
rect 32770 139200 32826 140000
rect 36818 139200 36874 140000
rect 40866 139200 40922 140000
rect 44914 139200 44970 140000
rect 48962 139200 49018 140000
rect 53010 139200 53066 140000
rect 57058 139200 57114 140000
rect 61106 139200 61162 140000
rect 65154 139200 65210 140000
rect 69202 139200 69258 140000
rect 73250 139200 73306 140000
rect 77298 139200 77354 140000
rect 81346 139200 81402 140000
rect 85394 139200 85450 140000
rect 89442 139200 89498 140000
rect 93490 139200 93546 140000
rect 97538 139200 97594 140000
rect 101586 139200 101642 140000
rect 105634 139200 105690 140000
rect 109682 139200 109738 140000
rect 113730 139200 113786 140000
rect 117778 139200 117834 140000
rect 121826 139200 121882 140000
rect 125874 139200 125930 140000
rect 129922 139200 129978 140000
rect 133970 139200 134026 140000
rect 138018 139200 138074 140000
rect 142066 139200 142122 140000
rect 146114 139200 146170 140000
rect 150162 139200 150218 140000
rect 154210 139200 154266 140000
rect 158258 139200 158314 140000
rect 162306 139200 162362 140000
rect 166354 139200 166410 140000
rect 170402 139200 170458 140000
rect 174450 139200 174506 140000
rect 178498 139200 178554 140000
rect 182546 139200 182602 140000
rect 186594 139200 186650 140000
rect 190642 139200 190698 140000
rect 194690 139200 194746 140000
rect 198738 139200 198794 140000
rect 202786 139200 202842 140000
rect 206834 139200 206890 140000
rect 210882 139200 210938 140000
rect 214930 139200 214986 140000
rect 218978 139200 219034 140000
rect 223026 139200 223082 140000
rect 227074 139200 227130 140000
rect 231122 139200 231178 140000
rect 235170 139200 235226 140000
rect 239218 139200 239274 140000
rect 243266 139200 243322 140000
rect 247314 139200 247370 140000
rect 251362 139200 251418 140000
rect 255410 139200 255466 140000
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16578 0 16634 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 40958 0 41014 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48778 0 48834 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57058 0 57114 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58438 0 58494 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61198 0 61254 800
rect 61658 0 61714 800
rect 62118 0 62174 800
rect 62578 0 62634 800
rect 63038 0 63094 800
rect 63498 0 63554 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64878 0 64934 800
rect 65338 0 65394 800
rect 65798 0 65854 800
rect 66258 0 66314 800
rect 66718 0 66774 800
rect 67178 0 67234 800
rect 67638 0 67694 800
rect 68098 0 68154 800
rect 68558 0 68614 800
rect 69018 0 69074 800
rect 69478 0 69534 800
rect 69938 0 69994 800
rect 70398 0 70454 800
rect 70858 0 70914 800
rect 71318 0 71374 800
rect 71778 0 71834 800
rect 72238 0 72294 800
rect 72698 0 72754 800
rect 73158 0 73214 800
rect 73618 0 73674 800
rect 74078 0 74134 800
rect 74538 0 74594 800
rect 74998 0 75054 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76378 0 76434 800
rect 76838 0 76894 800
rect 77298 0 77354 800
rect 77758 0 77814 800
rect 78218 0 78274 800
rect 78678 0 78734 800
rect 79138 0 79194 800
rect 79598 0 79654 800
rect 80058 0 80114 800
rect 80518 0 80574 800
rect 80978 0 81034 800
rect 81438 0 81494 800
rect 81898 0 81954 800
rect 82358 0 82414 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83738 0 83794 800
rect 84198 0 84254 800
rect 84658 0 84714 800
rect 85118 0 85174 800
rect 85578 0 85634 800
rect 86038 0 86094 800
rect 86498 0 86554 800
rect 86958 0 87014 800
rect 87418 0 87474 800
rect 87878 0 87934 800
rect 88338 0 88394 800
rect 88798 0 88854 800
rect 89258 0 89314 800
rect 89718 0 89774 800
rect 90178 0 90234 800
rect 90638 0 90694 800
rect 91098 0 91154 800
rect 91558 0 91614 800
rect 92018 0 92074 800
rect 92478 0 92534 800
rect 92938 0 92994 800
rect 93398 0 93454 800
rect 93858 0 93914 800
rect 94318 0 94374 800
rect 94778 0 94834 800
rect 95238 0 95294 800
rect 95698 0 95754 800
rect 96158 0 96214 800
rect 96618 0 96674 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 97998 0 98054 800
rect 98458 0 98514 800
rect 98918 0 98974 800
rect 99378 0 99434 800
rect 99838 0 99894 800
rect 100298 0 100354 800
rect 100758 0 100814 800
rect 101218 0 101274 800
rect 101678 0 101734 800
rect 102138 0 102194 800
rect 102598 0 102654 800
rect 103058 0 103114 800
rect 103518 0 103574 800
rect 103978 0 104034 800
rect 104438 0 104494 800
rect 104898 0 104954 800
rect 105358 0 105414 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 106738 0 106794 800
rect 107198 0 107254 800
rect 107658 0 107714 800
rect 108118 0 108174 800
rect 108578 0 108634 800
rect 109038 0 109094 800
rect 109498 0 109554 800
rect 109958 0 110014 800
rect 110418 0 110474 800
rect 110878 0 110934 800
rect 111338 0 111394 800
rect 111798 0 111854 800
rect 112258 0 112314 800
rect 112718 0 112774 800
rect 113178 0 113234 800
rect 113638 0 113694 800
rect 114098 0 114154 800
rect 114558 0 114614 800
rect 115018 0 115074 800
rect 115478 0 115534 800
rect 115938 0 115994 800
rect 116398 0 116454 800
rect 116858 0 116914 800
rect 117318 0 117374 800
rect 117778 0 117834 800
rect 118238 0 118294 800
rect 118698 0 118754 800
rect 119158 0 119214 800
rect 119618 0 119674 800
rect 120078 0 120134 800
rect 120538 0 120594 800
rect 120998 0 121054 800
rect 121458 0 121514 800
rect 121918 0 121974 800
rect 122378 0 122434 800
rect 122838 0 122894 800
rect 123298 0 123354 800
rect 123758 0 123814 800
rect 124218 0 124274 800
rect 124678 0 124734 800
rect 125138 0 125194 800
rect 125598 0 125654 800
rect 126058 0 126114 800
rect 126518 0 126574 800
rect 126978 0 127034 800
rect 127438 0 127494 800
rect 127898 0 127954 800
rect 128358 0 128414 800
rect 128818 0 128874 800
rect 129278 0 129334 800
rect 129738 0 129794 800
rect 130198 0 130254 800
rect 130658 0 130714 800
rect 131118 0 131174 800
rect 131578 0 131634 800
rect 132038 0 132094 800
rect 132498 0 132554 800
rect 132958 0 133014 800
rect 133418 0 133474 800
rect 133878 0 133934 800
rect 134338 0 134394 800
rect 134798 0 134854 800
rect 135258 0 135314 800
rect 135718 0 135774 800
rect 136178 0 136234 800
rect 136638 0 136694 800
rect 137098 0 137154 800
rect 137558 0 137614 800
rect 138018 0 138074 800
rect 138478 0 138534 800
rect 138938 0 138994 800
rect 139398 0 139454 800
rect 139858 0 139914 800
rect 140318 0 140374 800
rect 140778 0 140834 800
rect 141238 0 141294 800
rect 141698 0 141754 800
rect 142158 0 142214 800
rect 142618 0 142674 800
rect 143078 0 143134 800
rect 143538 0 143594 800
rect 143998 0 144054 800
rect 144458 0 144514 800
rect 144918 0 144974 800
rect 145378 0 145434 800
rect 145838 0 145894 800
rect 146298 0 146354 800
rect 146758 0 146814 800
rect 147218 0 147274 800
rect 147678 0 147734 800
rect 148138 0 148194 800
rect 148598 0 148654 800
rect 149058 0 149114 800
rect 149518 0 149574 800
rect 149978 0 150034 800
rect 150438 0 150494 800
rect 150898 0 150954 800
rect 151358 0 151414 800
rect 151818 0 151874 800
rect 152278 0 152334 800
rect 152738 0 152794 800
rect 153198 0 153254 800
rect 153658 0 153714 800
rect 154118 0 154174 800
rect 154578 0 154634 800
rect 155038 0 155094 800
rect 155498 0 155554 800
rect 155958 0 156014 800
rect 156418 0 156474 800
rect 156878 0 156934 800
rect 157338 0 157394 800
rect 157798 0 157854 800
rect 158258 0 158314 800
rect 158718 0 158774 800
rect 159178 0 159234 800
rect 159638 0 159694 800
rect 160098 0 160154 800
rect 160558 0 160614 800
rect 161018 0 161074 800
rect 161478 0 161534 800
rect 161938 0 161994 800
rect 162398 0 162454 800
rect 162858 0 162914 800
rect 163318 0 163374 800
rect 163778 0 163834 800
rect 164238 0 164294 800
rect 164698 0 164754 800
rect 165158 0 165214 800
rect 165618 0 165674 800
rect 166078 0 166134 800
rect 166538 0 166594 800
rect 166998 0 167054 800
rect 167458 0 167514 800
rect 167918 0 167974 800
rect 168378 0 168434 800
rect 168838 0 168894 800
rect 169298 0 169354 800
rect 169758 0 169814 800
rect 170218 0 170274 800
rect 170678 0 170734 800
rect 171138 0 171194 800
rect 171598 0 171654 800
rect 172058 0 172114 800
rect 172518 0 172574 800
rect 172978 0 173034 800
rect 173438 0 173494 800
rect 173898 0 173954 800
rect 174358 0 174414 800
rect 174818 0 174874 800
rect 175278 0 175334 800
rect 175738 0 175794 800
rect 176198 0 176254 800
rect 176658 0 176714 800
rect 177118 0 177174 800
rect 177578 0 177634 800
rect 178038 0 178094 800
rect 178498 0 178554 800
rect 178958 0 179014 800
rect 179418 0 179474 800
rect 179878 0 179934 800
rect 180338 0 180394 800
rect 180798 0 180854 800
rect 181258 0 181314 800
rect 181718 0 181774 800
rect 182178 0 182234 800
rect 182638 0 182694 800
rect 183098 0 183154 800
rect 183558 0 183614 800
rect 184018 0 184074 800
rect 184478 0 184534 800
rect 184938 0 184994 800
rect 185398 0 185454 800
rect 185858 0 185914 800
rect 186318 0 186374 800
rect 186778 0 186834 800
rect 187238 0 187294 800
rect 187698 0 187754 800
rect 188158 0 188214 800
rect 188618 0 188674 800
rect 189078 0 189134 800
rect 189538 0 189594 800
rect 189998 0 190054 800
rect 190458 0 190514 800
rect 190918 0 190974 800
rect 191378 0 191434 800
rect 191838 0 191894 800
rect 192298 0 192354 800
rect 192758 0 192814 800
rect 193218 0 193274 800
rect 193678 0 193734 800
rect 194138 0 194194 800
rect 194598 0 194654 800
rect 195058 0 195114 800
rect 195518 0 195574 800
rect 195978 0 196034 800
rect 196438 0 196494 800
rect 196898 0 196954 800
rect 197358 0 197414 800
rect 197818 0 197874 800
rect 198278 0 198334 800
rect 198738 0 198794 800
rect 199198 0 199254 800
rect 199658 0 199714 800
rect 200118 0 200174 800
rect 200578 0 200634 800
rect 201038 0 201094 800
rect 201498 0 201554 800
rect 201958 0 202014 800
rect 202418 0 202474 800
rect 202878 0 202934 800
rect 203338 0 203394 800
rect 203798 0 203854 800
rect 204258 0 204314 800
rect 204718 0 204774 800
rect 205178 0 205234 800
rect 205638 0 205694 800
rect 206098 0 206154 800
rect 206558 0 206614 800
rect 207018 0 207074 800
rect 207478 0 207534 800
rect 207938 0 207994 800
rect 208398 0 208454 800
rect 208858 0 208914 800
rect 209318 0 209374 800
rect 209778 0 209834 800
rect 210238 0 210294 800
rect 210698 0 210754 800
rect 211158 0 211214 800
rect 211618 0 211674 800
rect 212078 0 212134 800
rect 212538 0 212594 800
rect 212998 0 213054 800
rect 213458 0 213514 800
rect 213918 0 213974 800
rect 214378 0 214434 800
rect 214838 0 214894 800
rect 215298 0 215354 800
rect 215758 0 215814 800
rect 216218 0 216274 800
rect 216678 0 216734 800
rect 217138 0 217194 800
rect 217598 0 217654 800
rect 218058 0 218114 800
rect 218518 0 218574 800
rect 218978 0 219034 800
rect 219438 0 219494 800
rect 219898 0 219954 800
rect 220358 0 220414 800
rect 220818 0 220874 800
rect 221278 0 221334 800
rect 221738 0 221794 800
rect 222198 0 222254 800
rect 222658 0 222714 800
rect 223118 0 223174 800
rect 223578 0 223634 800
rect 224038 0 224094 800
rect 224498 0 224554 800
rect 224958 0 225014 800
rect 225418 0 225474 800
rect 225878 0 225934 800
rect 226338 0 226394 800
rect 226798 0 226854 800
rect 227258 0 227314 800
rect 227718 0 227774 800
rect 228178 0 228234 800
rect 228638 0 228694 800
rect 229098 0 229154 800
rect 229558 0 229614 800
rect 230018 0 230074 800
rect 230478 0 230534 800
rect 230938 0 230994 800
rect 231398 0 231454 800
rect 231858 0 231914 800
rect 232318 0 232374 800
rect 232778 0 232834 800
rect 233238 0 233294 800
rect 233698 0 233754 800
rect 234158 0 234214 800
rect 234618 0 234674 800
rect 235078 0 235134 800
rect 235538 0 235594 800
rect 235998 0 236054 800
rect 236458 0 236514 800
rect 236918 0 236974 800
rect 237378 0 237434 800
rect 237838 0 237894 800
rect 238298 0 238354 800
rect 238758 0 238814 800
rect 239218 0 239274 800
rect 239678 0 239734 800
rect 240138 0 240194 800
rect 240598 0 240654 800
rect 241058 0 241114 800
rect 241518 0 241574 800
rect 241978 0 242034 800
rect 242438 0 242494 800
rect 242898 0 242954 800
rect 243358 0 243414 800
rect 243818 0 243874 800
rect 244278 0 244334 800
rect 244738 0 244794 800
rect 245198 0 245254 800
rect 245658 0 245714 800
rect 246118 0 246174 800
rect 246578 0 246634 800
rect 247038 0 247094 800
rect 247498 0 247554 800
rect 247958 0 248014 800
rect 248418 0 248474 800
rect 248878 0 248934 800
rect 249338 0 249394 800
<< obsm2 >>
rect 938 139144 4378 139346
rect 4546 139144 8426 139346
rect 8594 139144 12474 139346
rect 12642 139144 16522 139346
rect 16690 139144 20570 139346
rect 20738 139144 24618 139346
rect 24786 139144 28666 139346
rect 28834 139144 32714 139346
rect 32882 139144 36762 139346
rect 36930 139144 40810 139346
rect 40978 139144 44858 139346
rect 45026 139144 48906 139346
rect 49074 139144 52954 139346
rect 53122 139144 57002 139346
rect 57170 139144 61050 139346
rect 61218 139144 65098 139346
rect 65266 139144 69146 139346
rect 69314 139144 73194 139346
rect 73362 139144 77242 139346
rect 77410 139144 81290 139346
rect 81458 139144 85338 139346
rect 85506 139144 89386 139346
rect 89554 139144 93434 139346
rect 93602 139144 97482 139346
rect 97650 139144 101530 139346
rect 101698 139144 105578 139346
rect 105746 139144 109626 139346
rect 109794 139144 113674 139346
rect 113842 139144 117722 139346
rect 117890 139144 121770 139346
rect 121938 139144 125818 139346
rect 125986 139144 129866 139346
rect 130034 139144 133914 139346
rect 134082 139144 137962 139346
rect 138130 139144 142010 139346
rect 142178 139144 146058 139346
rect 146226 139144 150106 139346
rect 150274 139144 154154 139346
rect 154322 139144 158202 139346
rect 158370 139144 162250 139346
rect 162418 139144 166298 139346
rect 166466 139144 170346 139346
rect 170514 139144 174394 139346
rect 174562 139144 178442 139346
rect 178610 139144 182490 139346
rect 182658 139144 186538 139346
rect 186706 139144 190586 139346
rect 190754 139144 194634 139346
rect 194802 139144 198682 139346
rect 198850 139144 202730 139346
rect 202898 139144 206778 139346
rect 206946 139144 210826 139346
rect 210994 139144 214874 139346
rect 215042 139144 218922 139346
rect 219090 139144 222970 139346
rect 223138 139144 227018 139346
rect 227186 139144 231066 139346
rect 231234 139144 235114 139346
rect 235282 139144 239162 139346
rect 239330 139144 243210 139346
rect 243378 139144 247258 139346
rect 247426 139144 251306 139346
rect 251474 139144 255354 139346
rect 255522 139144 255556 139346
rect 938 856 255556 139144
rect 938 734 10542 856
rect 10710 734 11002 856
rect 11170 734 11462 856
rect 11630 734 11922 856
rect 12090 734 12382 856
rect 12550 734 12842 856
rect 13010 734 13302 856
rect 13470 734 13762 856
rect 13930 734 14222 856
rect 14390 734 14682 856
rect 14850 734 15142 856
rect 15310 734 15602 856
rect 15770 734 16062 856
rect 16230 734 16522 856
rect 16690 734 16982 856
rect 17150 734 17442 856
rect 17610 734 17902 856
rect 18070 734 18362 856
rect 18530 734 18822 856
rect 18990 734 19282 856
rect 19450 734 19742 856
rect 19910 734 20202 856
rect 20370 734 20662 856
rect 20830 734 21122 856
rect 21290 734 21582 856
rect 21750 734 22042 856
rect 22210 734 22502 856
rect 22670 734 22962 856
rect 23130 734 23422 856
rect 23590 734 23882 856
rect 24050 734 24342 856
rect 24510 734 24802 856
rect 24970 734 25262 856
rect 25430 734 25722 856
rect 25890 734 26182 856
rect 26350 734 26642 856
rect 26810 734 27102 856
rect 27270 734 27562 856
rect 27730 734 28022 856
rect 28190 734 28482 856
rect 28650 734 28942 856
rect 29110 734 29402 856
rect 29570 734 29862 856
rect 30030 734 30322 856
rect 30490 734 30782 856
rect 30950 734 31242 856
rect 31410 734 31702 856
rect 31870 734 32162 856
rect 32330 734 32622 856
rect 32790 734 33082 856
rect 33250 734 33542 856
rect 33710 734 34002 856
rect 34170 734 34462 856
rect 34630 734 34922 856
rect 35090 734 35382 856
rect 35550 734 35842 856
rect 36010 734 36302 856
rect 36470 734 36762 856
rect 36930 734 37222 856
rect 37390 734 37682 856
rect 37850 734 38142 856
rect 38310 734 38602 856
rect 38770 734 39062 856
rect 39230 734 39522 856
rect 39690 734 39982 856
rect 40150 734 40442 856
rect 40610 734 40902 856
rect 41070 734 41362 856
rect 41530 734 41822 856
rect 41990 734 42282 856
rect 42450 734 42742 856
rect 42910 734 43202 856
rect 43370 734 43662 856
rect 43830 734 44122 856
rect 44290 734 44582 856
rect 44750 734 45042 856
rect 45210 734 45502 856
rect 45670 734 45962 856
rect 46130 734 46422 856
rect 46590 734 46882 856
rect 47050 734 47342 856
rect 47510 734 47802 856
rect 47970 734 48262 856
rect 48430 734 48722 856
rect 48890 734 49182 856
rect 49350 734 49642 856
rect 49810 734 50102 856
rect 50270 734 50562 856
rect 50730 734 51022 856
rect 51190 734 51482 856
rect 51650 734 51942 856
rect 52110 734 52402 856
rect 52570 734 52862 856
rect 53030 734 53322 856
rect 53490 734 53782 856
rect 53950 734 54242 856
rect 54410 734 54702 856
rect 54870 734 55162 856
rect 55330 734 55622 856
rect 55790 734 56082 856
rect 56250 734 56542 856
rect 56710 734 57002 856
rect 57170 734 57462 856
rect 57630 734 57922 856
rect 58090 734 58382 856
rect 58550 734 58842 856
rect 59010 734 59302 856
rect 59470 734 59762 856
rect 59930 734 60222 856
rect 60390 734 60682 856
rect 60850 734 61142 856
rect 61310 734 61602 856
rect 61770 734 62062 856
rect 62230 734 62522 856
rect 62690 734 62982 856
rect 63150 734 63442 856
rect 63610 734 63902 856
rect 64070 734 64362 856
rect 64530 734 64822 856
rect 64990 734 65282 856
rect 65450 734 65742 856
rect 65910 734 66202 856
rect 66370 734 66662 856
rect 66830 734 67122 856
rect 67290 734 67582 856
rect 67750 734 68042 856
rect 68210 734 68502 856
rect 68670 734 68962 856
rect 69130 734 69422 856
rect 69590 734 69882 856
rect 70050 734 70342 856
rect 70510 734 70802 856
rect 70970 734 71262 856
rect 71430 734 71722 856
rect 71890 734 72182 856
rect 72350 734 72642 856
rect 72810 734 73102 856
rect 73270 734 73562 856
rect 73730 734 74022 856
rect 74190 734 74482 856
rect 74650 734 74942 856
rect 75110 734 75402 856
rect 75570 734 75862 856
rect 76030 734 76322 856
rect 76490 734 76782 856
rect 76950 734 77242 856
rect 77410 734 77702 856
rect 77870 734 78162 856
rect 78330 734 78622 856
rect 78790 734 79082 856
rect 79250 734 79542 856
rect 79710 734 80002 856
rect 80170 734 80462 856
rect 80630 734 80922 856
rect 81090 734 81382 856
rect 81550 734 81842 856
rect 82010 734 82302 856
rect 82470 734 82762 856
rect 82930 734 83222 856
rect 83390 734 83682 856
rect 83850 734 84142 856
rect 84310 734 84602 856
rect 84770 734 85062 856
rect 85230 734 85522 856
rect 85690 734 85982 856
rect 86150 734 86442 856
rect 86610 734 86902 856
rect 87070 734 87362 856
rect 87530 734 87822 856
rect 87990 734 88282 856
rect 88450 734 88742 856
rect 88910 734 89202 856
rect 89370 734 89662 856
rect 89830 734 90122 856
rect 90290 734 90582 856
rect 90750 734 91042 856
rect 91210 734 91502 856
rect 91670 734 91962 856
rect 92130 734 92422 856
rect 92590 734 92882 856
rect 93050 734 93342 856
rect 93510 734 93802 856
rect 93970 734 94262 856
rect 94430 734 94722 856
rect 94890 734 95182 856
rect 95350 734 95642 856
rect 95810 734 96102 856
rect 96270 734 96562 856
rect 96730 734 97022 856
rect 97190 734 97482 856
rect 97650 734 97942 856
rect 98110 734 98402 856
rect 98570 734 98862 856
rect 99030 734 99322 856
rect 99490 734 99782 856
rect 99950 734 100242 856
rect 100410 734 100702 856
rect 100870 734 101162 856
rect 101330 734 101622 856
rect 101790 734 102082 856
rect 102250 734 102542 856
rect 102710 734 103002 856
rect 103170 734 103462 856
rect 103630 734 103922 856
rect 104090 734 104382 856
rect 104550 734 104842 856
rect 105010 734 105302 856
rect 105470 734 105762 856
rect 105930 734 106222 856
rect 106390 734 106682 856
rect 106850 734 107142 856
rect 107310 734 107602 856
rect 107770 734 108062 856
rect 108230 734 108522 856
rect 108690 734 108982 856
rect 109150 734 109442 856
rect 109610 734 109902 856
rect 110070 734 110362 856
rect 110530 734 110822 856
rect 110990 734 111282 856
rect 111450 734 111742 856
rect 111910 734 112202 856
rect 112370 734 112662 856
rect 112830 734 113122 856
rect 113290 734 113582 856
rect 113750 734 114042 856
rect 114210 734 114502 856
rect 114670 734 114962 856
rect 115130 734 115422 856
rect 115590 734 115882 856
rect 116050 734 116342 856
rect 116510 734 116802 856
rect 116970 734 117262 856
rect 117430 734 117722 856
rect 117890 734 118182 856
rect 118350 734 118642 856
rect 118810 734 119102 856
rect 119270 734 119562 856
rect 119730 734 120022 856
rect 120190 734 120482 856
rect 120650 734 120942 856
rect 121110 734 121402 856
rect 121570 734 121862 856
rect 122030 734 122322 856
rect 122490 734 122782 856
rect 122950 734 123242 856
rect 123410 734 123702 856
rect 123870 734 124162 856
rect 124330 734 124622 856
rect 124790 734 125082 856
rect 125250 734 125542 856
rect 125710 734 126002 856
rect 126170 734 126462 856
rect 126630 734 126922 856
rect 127090 734 127382 856
rect 127550 734 127842 856
rect 128010 734 128302 856
rect 128470 734 128762 856
rect 128930 734 129222 856
rect 129390 734 129682 856
rect 129850 734 130142 856
rect 130310 734 130602 856
rect 130770 734 131062 856
rect 131230 734 131522 856
rect 131690 734 131982 856
rect 132150 734 132442 856
rect 132610 734 132902 856
rect 133070 734 133362 856
rect 133530 734 133822 856
rect 133990 734 134282 856
rect 134450 734 134742 856
rect 134910 734 135202 856
rect 135370 734 135662 856
rect 135830 734 136122 856
rect 136290 734 136582 856
rect 136750 734 137042 856
rect 137210 734 137502 856
rect 137670 734 137962 856
rect 138130 734 138422 856
rect 138590 734 138882 856
rect 139050 734 139342 856
rect 139510 734 139802 856
rect 139970 734 140262 856
rect 140430 734 140722 856
rect 140890 734 141182 856
rect 141350 734 141642 856
rect 141810 734 142102 856
rect 142270 734 142562 856
rect 142730 734 143022 856
rect 143190 734 143482 856
rect 143650 734 143942 856
rect 144110 734 144402 856
rect 144570 734 144862 856
rect 145030 734 145322 856
rect 145490 734 145782 856
rect 145950 734 146242 856
rect 146410 734 146702 856
rect 146870 734 147162 856
rect 147330 734 147622 856
rect 147790 734 148082 856
rect 148250 734 148542 856
rect 148710 734 149002 856
rect 149170 734 149462 856
rect 149630 734 149922 856
rect 150090 734 150382 856
rect 150550 734 150842 856
rect 151010 734 151302 856
rect 151470 734 151762 856
rect 151930 734 152222 856
rect 152390 734 152682 856
rect 152850 734 153142 856
rect 153310 734 153602 856
rect 153770 734 154062 856
rect 154230 734 154522 856
rect 154690 734 154982 856
rect 155150 734 155442 856
rect 155610 734 155902 856
rect 156070 734 156362 856
rect 156530 734 156822 856
rect 156990 734 157282 856
rect 157450 734 157742 856
rect 157910 734 158202 856
rect 158370 734 158662 856
rect 158830 734 159122 856
rect 159290 734 159582 856
rect 159750 734 160042 856
rect 160210 734 160502 856
rect 160670 734 160962 856
rect 161130 734 161422 856
rect 161590 734 161882 856
rect 162050 734 162342 856
rect 162510 734 162802 856
rect 162970 734 163262 856
rect 163430 734 163722 856
rect 163890 734 164182 856
rect 164350 734 164642 856
rect 164810 734 165102 856
rect 165270 734 165562 856
rect 165730 734 166022 856
rect 166190 734 166482 856
rect 166650 734 166942 856
rect 167110 734 167402 856
rect 167570 734 167862 856
rect 168030 734 168322 856
rect 168490 734 168782 856
rect 168950 734 169242 856
rect 169410 734 169702 856
rect 169870 734 170162 856
rect 170330 734 170622 856
rect 170790 734 171082 856
rect 171250 734 171542 856
rect 171710 734 172002 856
rect 172170 734 172462 856
rect 172630 734 172922 856
rect 173090 734 173382 856
rect 173550 734 173842 856
rect 174010 734 174302 856
rect 174470 734 174762 856
rect 174930 734 175222 856
rect 175390 734 175682 856
rect 175850 734 176142 856
rect 176310 734 176602 856
rect 176770 734 177062 856
rect 177230 734 177522 856
rect 177690 734 177982 856
rect 178150 734 178442 856
rect 178610 734 178902 856
rect 179070 734 179362 856
rect 179530 734 179822 856
rect 179990 734 180282 856
rect 180450 734 180742 856
rect 180910 734 181202 856
rect 181370 734 181662 856
rect 181830 734 182122 856
rect 182290 734 182582 856
rect 182750 734 183042 856
rect 183210 734 183502 856
rect 183670 734 183962 856
rect 184130 734 184422 856
rect 184590 734 184882 856
rect 185050 734 185342 856
rect 185510 734 185802 856
rect 185970 734 186262 856
rect 186430 734 186722 856
rect 186890 734 187182 856
rect 187350 734 187642 856
rect 187810 734 188102 856
rect 188270 734 188562 856
rect 188730 734 189022 856
rect 189190 734 189482 856
rect 189650 734 189942 856
rect 190110 734 190402 856
rect 190570 734 190862 856
rect 191030 734 191322 856
rect 191490 734 191782 856
rect 191950 734 192242 856
rect 192410 734 192702 856
rect 192870 734 193162 856
rect 193330 734 193622 856
rect 193790 734 194082 856
rect 194250 734 194542 856
rect 194710 734 195002 856
rect 195170 734 195462 856
rect 195630 734 195922 856
rect 196090 734 196382 856
rect 196550 734 196842 856
rect 197010 734 197302 856
rect 197470 734 197762 856
rect 197930 734 198222 856
rect 198390 734 198682 856
rect 198850 734 199142 856
rect 199310 734 199602 856
rect 199770 734 200062 856
rect 200230 734 200522 856
rect 200690 734 200982 856
rect 201150 734 201442 856
rect 201610 734 201902 856
rect 202070 734 202362 856
rect 202530 734 202822 856
rect 202990 734 203282 856
rect 203450 734 203742 856
rect 203910 734 204202 856
rect 204370 734 204662 856
rect 204830 734 205122 856
rect 205290 734 205582 856
rect 205750 734 206042 856
rect 206210 734 206502 856
rect 206670 734 206962 856
rect 207130 734 207422 856
rect 207590 734 207882 856
rect 208050 734 208342 856
rect 208510 734 208802 856
rect 208970 734 209262 856
rect 209430 734 209722 856
rect 209890 734 210182 856
rect 210350 734 210642 856
rect 210810 734 211102 856
rect 211270 734 211562 856
rect 211730 734 212022 856
rect 212190 734 212482 856
rect 212650 734 212942 856
rect 213110 734 213402 856
rect 213570 734 213862 856
rect 214030 734 214322 856
rect 214490 734 214782 856
rect 214950 734 215242 856
rect 215410 734 215702 856
rect 215870 734 216162 856
rect 216330 734 216622 856
rect 216790 734 217082 856
rect 217250 734 217542 856
rect 217710 734 218002 856
rect 218170 734 218462 856
rect 218630 734 218922 856
rect 219090 734 219382 856
rect 219550 734 219842 856
rect 220010 734 220302 856
rect 220470 734 220762 856
rect 220930 734 221222 856
rect 221390 734 221682 856
rect 221850 734 222142 856
rect 222310 734 222602 856
rect 222770 734 223062 856
rect 223230 734 223522 856
rect 223690 734 223982 856
rect 224150 734 224442 856
rect 224610 734 224902 856
rect 225070 734 225362 856
rect 225530 734 225822 856
rect 225990 734 226282 856
rect 226450 734 226742 856
rect 226910 734 227202 856
rect 227370 734 227662 856
rect 227830 734 228122 856
rect 228290 734 228582 856
rect 228750 734 229042 856
rect 229210 734 229502 856
rect 229670 734 229962 856
rect 230130 734 230422 856
rect 230590 734 230882 856
rect 231050 734 231342 856
rect 231510 734 231802 856
rect 231970 734 232262 856
rect 232430 734 232722 856
rect 232890 734 233182 856
rect 233350 734 233642 856
rect 233810 734 234102 856
rect 234270 734 234562 856
rect 234730 734 235022 856
rect 235190 734 235482 856
rect 235650 734 235942 856
rect 236110 734 236402 856
rect 236570 734 236862 856
rect 237030 734 237322 856
rect 237490 734 237782 856
rect 237950 734 238242 856
rect 238410 734 238702 856
rect 238870 734 239162 856
rect 239330 734 239622 856
rect 239790 734 240082 856
rect 240250 734 240542 856
rect 240710 734 241002 856
rect 241170 734 241462 856
rect 241630 734 241922 856
rect 242090 734 242382 856
rect 242550 734 242842 856
rect 243010 734 243302 856
rect 243470 734 243762 856
rect 243930 734 244222 856
rect 244390 734 244682 856
rect 244850 734 245142 856
rect 245310 734 245602 856
rect 245770 734 246062 856
rect 246230 734 246522 856
rect 246690 734 246982 856
rect 247150 734 247442 856
rect 247610 734 247902 856
rect 248070 734 248362 856
rect 248530 734 248822 856
rect 248990 734 249282 856
rect 249450 734 255556 856
<< metal3 >>
rect 0 134648 800 134768
rect 0 132200 800 132320
rect 0 129752 800 129872
rect 0 127304 800 127424
rect 0 124856 800 124976
rect 0 122408 800 122528
rect 0 119960 800 120080
rect 0 117512 800 117632
rect 0 115064 800 115184
rect 0 112616 800 112736
rect 0 110168 800 110288
rect 0 107720 800 107840
rect 0 105272 800 105392
rect 0 102824 800 102944
rect 0 100376 800 100496
rect 0 97928 800 98048
rect 0 95480 800 95600
rect 0 93032 800 93152
rect 0 90584 800 90704
rect 0 88136 800 88256
rect 0 85688 800 85808
rect 0 83240 800 83360
rect 0 80792 800 80912
rect 0 78344 800 78464
rect 0 75896 800 76016
rect 0 73448 800 73568
rect 0 71000 800 71120
rect 0 68552 800 68672
rect 0 66104 800 66224
rect 0 63656 800 63776
rect 0 61208 800 61328
rect 0 58760 800 58880
rect 0 56312 800 56432
rect 0 53864 800 53984
rect 0 51416 800 51536
rect 0 48968 800 49088
rect 0 46520 800 46640
rect 0 44072 800 44192
rect 0 41624 800 41744
rect 0 39176 800 39296
rect 0 36728 800 36848
rect 0 34280 800 34400
rect 0 31832 800 31952
rect 0 29384 800 29504
rect 0 26936 800 27056
rect 0 24488 800 24608
rect 0 22040 800 22160
rect 0 19592 800 19712
rect 0 17144 800 17264
rect 0 14696 800 14816
rect 0 12248 800 12368
rect 0 9800 800 9920
rect 0 7352 800 7472
rect 0 4904 800 5024
<< obsm3 >>
rect 798 134848 250286 137665
rect 880 134568 250286 134848
rect 798 132400 250286 134568
rect 880 132120 250286 132400
rect 798 129952 250286 132120
rect 880 129672 250286 129952
rect 798 127504 250286 129672
rect 880 127224 250286 127504
rect 798 125056 250286 127224
rect 880 124776 250286 125056
rect 798 122608 250286 124776
rect 880 122328 250286 122608
rect 798 120160 250286 122328
rect 880 119880 250286 120160
rect 798 117712 250286 119880
rect 880 117432 250286 117712
rect 798 115264 250286 117432
rect 880 114984 250286 115264
rect 798 112816 250286 114984
rect 880 112536 250286 112816
rect 798 110368 250286 112536
rect 880 110088 250286 110368
rect 798 107920 250286 110088
rect 880 107640 250286 107920
rect 798 105472 250286 107640
rect 880 105192 250286 105472
rect 798 103024 250286 105192
rect 880 102744 250286 103024
rect 798 100576 250286 102744
rect 880 100296 250286 100576
rect 798 98128 250286 100296
rect 880 97848 250286 98128
rect 798 95680 250286 97848
rect 880 95400 250286 95680
rect 798 93232 250286 95400
rect 880 92952 250286 93232
rect 798 90784 250286 92952
rect 880 90504 250286 90784
rect 798 88336 250286 90504
rect 880 88056 250286 88336
rect 798 85888 250286 88056
rect 880 85608 250286 85888
rect 798 83440 250286 85608
rect 880 83160 250286 83440
rect 798 80992 250286 83160
rect 880 80712 250286 80992
rect 798 78544 250286 80712
rect 880 78264 250286 78544
rect 798 76096 250286 78264
rect 880 75816 250286 76096
rect 798 73648 250286 75816
rect 880 73368 250286 73648
rect 798 71200 250286 73368
rect 880 70920 250286 71200
rect 798 68752 250286 70920
rect 880 68472 250286 68752
rect 798 66304 250286 68472
rect 880 66024 250286 66304
rect 798 63856 250286 66024
rect 880 63576 250286 63856
rect 798 61408 250286 63576
rect 880 61128 250286 61408
rect 798 58960 250286 61128
rect 880 58680 250286 58960
rect 798 56512 250286 58680
rect 880 56232 250286 56512
rect 798 54064 250286 56232
rect 880 53784 250286 54064
rect 798 51616 250286 53784
rect 880 51336 250286 51616
rect 798 49168 250286 51336
rect 880 48888 250286 49168
rect 798 46720 250286 48888
rect 880 46440 250286 46720
rect 798 44272 250286 46440
rect 880 43992 250286 44272
rect 798 41824 250286 43992
rect 880 41544 250286 41824
rect 798 39376 250286 41544
rect 880 39096 250286 39376
rect 798 36928 250286 39096
rect 880 36648 250286 36928
rect 798 34480 250286 36648
rect 880 34200 250286 34480
rect 798 32032 250286 34200
rect 880 31752 250286 32032
rect 798 29584 250286 31752
rect 880 29304 250286 29584
rect 798 27136 250286 29304
rect 880 26856 250286 27136
rect 798 24688 250286 26856
rect 880 24408 250286 24688
rect 798 22240 250286 24408
rect 880 21960 250286 22240
rect 798 19792 250286 21960
rect 880 19512 250286 19792
rect 798 17344 250286 19512
rect 880 17064 250286 17344
rect 798 14896 250286 17064
rect 880 14616 250286 14896
rect 798 12448 250286 14616
rect 880 12168 250286 12448
rect 798 10000 250286 12168
rect 880 9720 250286 10000
rect 798 7552 250286 9720
rect 880 7272 250286 7552
rect 798 5104 250286 7272
rect 880 4824 250286 5104
rect 798 2143 250286 4824
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
rect 142448 2128 142768 137680
rect 157808 2128 158128 137680
rect 173168 2128 173488 137680
rect 188528 2128 188848 137680
rect 203888 2128 204208 137680
rect 219248 2128 219568 137680
rect 234608 2128 234928 137680
rect 249968 2128 250288 137680
<< labels >>
rlabel metal2 s 245658 0 245714 800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 146114 139200 146170 140000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 162306 139200 162362 140000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 178498 139200 178554 140000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 194690 139200 194746 140000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 210882 139200 210938 140000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 227074 139200 227130 140000 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 243266 139200 243322 140000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 4904 800 5024 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 14696 800 14816 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 24488 800 24608 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 247498 0 247554 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 34280 800 34400 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 44072 800 44192 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 53864 800 53984 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 63656 800 63776 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 73448 800 73568 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 83240 800 83360 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 93032 800 93152 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 102824 800 102944 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 112616 800 112736 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal2 s 16578 139200 16634 140000 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal2 s 32770 139200 32826 140000 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 48962 139200 49018 140000 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal2 s 65154 139200 65210 140000 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 81346 139200 81402 140000 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 97538 139200 97594 140000 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 113730 139200 113786 140000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 129922 139200 129978 140000 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 235998 0 236054 800 6 io_in[0]
port 30 nsew signal input
rlabel metal2 s 36818 139200 36874 140000 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 53010 139200 53066 140000 6 io_in[11]
port 32 nsew signal input
rlabel metal2 s 69202 139200 69258 140000 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 85394 139200 85450 140000 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 101586 139200 101642 140000 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 117778 139200 117834 140000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 133970 139200 134026 140000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 150162 139200 150218 140000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 166354 139200 166410 140000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 182546 139200 182602 140000 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 198738 139200 198794 140000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 214930 139200 214986 140000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 231122 139200 231178 140000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 247314 139200 247370 140000 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 240138 0 240194 800 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 241518 0 241574 800 6 io_in[4]
port 62 nsew signal input
rlabel metal2 s 242898 0 242954 800 6 io_in[5]
port 63 nsew signal input
rlabel metal2 s 244278 0 244334 800 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 4434 139200 4490 140000 6 io_in[8]
port 66 nsew signal input
rlabel metal2 s 20626 139200 20682 140000 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 44914 139200 44970 140000 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 61106 139200 61162 140000 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 77298 139200 77354 140000 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 93490 139200 93546 140000 6 io_oeb[13]
port 72 nsew signal output
rlabel metal2 s 109682 139200 109738 140000 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 125874 139200 125930 140000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 142066 139200 142122 140000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 158258 139200 158314 140000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 174450 139200 174506 140000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 190642 139200 190698 140000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 238298 0 238354 800 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 206834 139200 206890 140000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 223026 139200 223082 140000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 239218 139200 239274 140000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 255410 139200 255466 140000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 239678 0 239734 800 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 100376 800 100496 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 119960 800 120080 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 io_oeb[3]
port 99 nsew signal output
rlabel metal2 s 242438 0 242494 800 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 243818 0 243874 800 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 245198 0 245254 800 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 247038 0 247094 800 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 12530 139200 12586 140000 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 28722 139200 28778 140000 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 io_out[0]
port 106 nsew signal output
rlabel metal2 s 40866 139200 40922 140000 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 57058 139200 57114 140000 6 io_out[11]
port 108 nsew signal output
rlabel metal2 s 73250 139200 73306 140000 6 io_out[12]
port 109 nsew signal output
rlabel metal2 s 89442 139200 89498 140000 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 105634 139200 105690 140000 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 121826 139200 121882 140000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 138018 139200 138074 140000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 154210 139200 154266 140000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 170402 139200 170458 140000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 186594 139200 186650 140000 6 io_out[19]
port 116 nsew signal output
rlabel metal2 s 237838 0 237894 800 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 202786 139200 202842 140000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 218978 139200 219034 140000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 235170 139200 235226 140000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 251362 139200 251418 140000 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 132200 800 132320 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 240598 0 240654 800 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 241978 0 242034 800 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 243358 0 243414 800 6 io_out[5]
port 139 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 246578 0 246634 800 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 8482 139200 8538 140000 6 io_out[8]
port 142 nsew signal output
rlabel metal2 s 24674 139200 24730 140000 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 167918 0 167974 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 168838 0 168894 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 172978 0 173034 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 175278 0 175334 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 176658 0 176714 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 143078 0 143134 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 149978 0 150034 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 155038 0 155094 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 158258 0 158314 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 160558 0 160614 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 162398 0 162454 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 163778 0 163834 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 177118 0 177174 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 224038 0 224094 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 224498 0 224554 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 224958 0 225014 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 225878 0 225934 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 229098 0 229154 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 229558 0 229614 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 182178 0 182234 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 233698 0 233754 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 234158 0 234214 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 234618 0 234674 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 235538 0 235594 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 190918 0 190974 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 191838 0 191894 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 192298 0 192354 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 197818 0 197874 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 198738 0 198794 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 200578 0 200634 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 202418 0 202474 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 204258 0 204314 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 205178 0 205234 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 207938 0 207994 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 210698 0 210754 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 211158 0 211214 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 216218 0 216274 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 216678 0 216734 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 217598 0 217654 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 218518 0 218574 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 221278 0 221334 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 248418 0 248474 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 249338 0 249394 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 137680 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 137680 6 vssd1
port 533 nsew ground bidirectional
rlabel metal2 s 10598 0 10654 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 260000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9663686
string GDS_FILE /root/eda/caravel_user_project/openlane/TOP_digital/runs/23_10_15_15_48/results/signoff/TOP_digital.magic.gds
string GDS_START 100956
<< end >>

